`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/19/2021 04:32:14 PM
// Design Name: 
// Module Name: addressgen_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module addressgen_unit(
    input  [`DataBusBits-1:0] reg1,
    input  [`DataBusBits-1:0] instruction,
    output reg [`DataBusBits-1:0] address
    );
    
    
endmodule
